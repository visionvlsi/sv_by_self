interface counter_intf;

logic clk,rst;
logic ld, ud;
logic [15:0]loadin;
logic [15:0]count;

endinterface