interface aif();
  logic [3:0]a,b;
  logic [7:0]prod;
endinterface