class transaction;

rand bit rst, ld, ud;
rand bit [15:0]loadin;
bit clk;
bit [15:0]count;
endclass