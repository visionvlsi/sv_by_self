//////////////////////////	Interface
 
interface mux_intf();
logic y;
logic [3:0]i;
logic [1:0]s;
endinterface
