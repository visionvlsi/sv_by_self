/////////////////////////////////	Transaction class

class transaction;
randc bit [3:0] i;
randc bit [1:0] s;
bit  y;
endclass
