`include "counter16.sv"
`include "tran.sv"
`include "gen.sv"
`include "intf.sv"
`include "drvr.sv"
`include "mon.sv"
//`include "sco.sv"
`include "env.sv"
`include "tb.sv"