`include "adder.sv"
`include "trans.sv"
`include "gen.sv"
`include "intf.sv"
`include "drv.sv"
`include "moni.sv"
`include "sco.sv"
`include "env.sv"
`include "test.sv"
`include "tb_top.sv"