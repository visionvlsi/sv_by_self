interface adder_intf;

logic [7:0]a,b;
logic [8:0]sum;

endinterface