interface intf();
  
  logic [7:0]a,b;
  logic enable;
  logic [3:0]command;
  logic [15:0]out;
  
  endinterface