//Design 4-bit adder

module mult(a,b,prod);
input [3:0]a,b;
output [7:0]prod;
assign prod=a*b;
endmodule

